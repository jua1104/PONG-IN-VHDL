LIBRARY ieee;
USE ieee.std_logic_1164.all;
-----------------------------------------------------------------
ENTITY PRINT_SCORE IS
PORT( binM : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		sseg : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		sseg_2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
);
END ENTITY PRINT_SCORE;
-------------------------------------------------------------------
ARCHITECTURE behaviour OF PRINT_SCORE IS
SIGNAL sseg_ou : STD_LOGIC_VECTOR(13 DOWNTO 0);
BEGIN
--sseg_ou <= sseg & sseg_2;
sseg <= sseg_ou(13 DOWNTO 7);
sseg_2 <= sseg_ou(6 DOWNTO 0);
WITH binM SELECT
sseg_ou<=
"10000001000000" WHEN "00000000", -- 00
"10000001111001" WHEN "00000001", -- 01
"10000000100100" WHEN "00000010", -- 02
"10000000110000" WHEN "00000011", -- 03
"10000000011001" WHEN "00000100", -- 04
"10000000010010" WHEN "00000101", -- 05
"10000000000010" WHEN "00000110", -- 06
"10000001111000" WHEN "00000111", -- 07
"10000000000000" WHEN "00001000", -- 08
"10000000010000" WHEN "00001001", -- 09
"11110011000000" WHEN "00001010", -- 10
"11110011111001" WHEN "00001011", -- 11
"11110010100100" WHEN "00001100", -- 12
"11110010110000" WHEN "00001101", -- 13
"11110010011001" WHEN "00001110", -- 14
"11110010010010" WHEN "00001111", -- 15
"11110010000010" WHEN "00010000", -- 16
"11110011111000" WHEN "00010001", -- 17
"11110010000000" WHEN "00010010", -- 18
"11110010010000" WHEN "00010011", -- 19
"01001001000000" WHEN "00010100", -- 20
"01001001111001" WHEN "00010101", -- 21
"01001000100100" WHEN "00010110", -- 22
"01001000110000" WHEN "00010111", -- 23
"01001000011001" WHEN "00011000", -- 24
"01001000010010" WHEN "00011001", -- 25
"01001000000010" WHEN "00011010", -- 26
"01001001111000" WHEN "00011011", -- 27
"01001000000000" WHEN "00011100", -- 28
"01001000010000" WHEN "00011101", -- 29
"01100001000000" WHEN "00011110", -- 30
"01100001111001" WHEN "00011111", -- 31
"01100000100100" WHEN "00100000", -- 32
"01100000110000" WHEN "00100001", -- 33
"01100000011001" WHEN "00100010", -- 34
"01100000010010" WHEN "00100011", -- 35
"01100000000010" WHEN "00100100", -- 36
"01100001111000" WHEN "00100101", -- 37
"01100000000000" WHEN "00100110", -- 38
"01100000010000" WHEN "00100111", -- 39
"00110011000000" WHEN "00101000", -- 40
"00110011111001" WHEN "00101001", -- 41
"00110010100100" WHEN "00101010", -- 42
"00110010110000" WHEN "00101011", -- 43
"00110010011001" WHEN "00101100", -- 44
"00110010010010" WHEN "00101101", -- 45
"00110010000010" WHEN "00101110", -- 46
"00110011111000" WHEN "00101111", -- 47
"00110010000000" WHEN "00110000", -- 48
"00110010010000" WHEN "00110001", -- 49
"00100101000000" WHEN "00110010", -- 50
"00100101111001" WHEN "00110011", -- 51
"00100100100100" WHEN "00110100", -- 52
"00100100110000" WHEN "00110101", -- 53
"00100100011001" WHEN "00110110", -- 54
"00100100010010" WHEN "00110111", -- 55
"00100100000010" WHEN "00111000", -- 56
"00100101111000" WHEN "00111001", -- 57
"00100100000000" WHEN "00111010", -- 58
"00100100010000" WHEN "00111011", -- 59
"00000101000000" WHEN "00111100", -- 60
"00000101111001" WHEN "00111101", -- 61
"00000100100100" WHEN "00111110", -- 62
"00000100110000" WHEN "00111111", -- 63
"00000100011001" WHEN "01000000", -- 64
"00000100010010" WHEN "01000001", -- 65
"00000100000010" WHEN "01000010", -- 66
"00000101111000" WHEN "01000011", -- 67
"00000100000000" WHEN "01000100", -- 68
"00000100010000" WHEN "01000101", -- 69
"11110001000000" WHEN "01000110", -- 70
"11110001111001" WHEN "01000111", -- 71
"11110000100100" WHEN "01001000", -- 72
"11110000110000" WHEN "01001001", -- 73
"11110000011001" WHEN "01001010", -- 74
"11110000010010" WHEN "01001011", -- 75
"11110000000010" WHEN "01001100", -- 76
"11110001111000" WHEN "01001101", -- 77
"11110000000000" WHEN "01001110", -- 78
"11110000010000" WHEN "01001111", -- 79
"00000001000000" WHEN "01010000", -- 80
"00000001111001" WHEN "01010001", -- 81
"00000000000000" WHEN OTHERS;
END behaviour;